module sipo_reg_tb;



endmodule
