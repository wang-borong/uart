module baud_gen (
    input sys_clk,
    input rst_n,
    output baud_clk
);


endmodule
