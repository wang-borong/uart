module parity_chk_tb;




endmodule
